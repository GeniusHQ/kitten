module main

pub enum Platform {
	unknown = -1
	any
	discord
	guilded
}