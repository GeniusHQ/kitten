module discord

pub type Snowflake = string