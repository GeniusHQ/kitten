module universe

pub enum Platform as int {
	unknown = -1
	any
	discord
	guilded
}