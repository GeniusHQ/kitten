module gateway

type Snowflake = string