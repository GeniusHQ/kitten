module gateway

struct GatewayBotResponse {
	url    string
	shards int
	// Todo: add session_start_limit
}
